module sprite_rom (
  input   [9:0]   addr_i,
  output  [63:0]  data_o
);

  localparam int AddrWidth = 10;
  localparam int DataWidth = 64;

  localparam logic [0:2**AddrWidth-1][DataWidth-1:0] ROM = {
    // code x00
    64'h0000000100000000,
    64'h0000000100000000,
    64'h0000000100000000,
    64'h0000001110000000,
    64'h0000001110000000,
    64'h0002001110020000,
    64'h0002001110020000,
    64'h0001011111010000,
    64'h2001711211710020,
    64'h2007112221170020,
    64'h1001112121110010,
    64'h1011111111111010,
    64'h1111121112111110,
    64'h1110221112201110,
    64'h1100220102200110,
    64'h1000000100000010,
    // code x01
    64'h0000001000000000,
    64'h0000001000000000,
    64'h0000001000000000,
    64'h0000011100000000,
    64'h0000011100200000,
    64'h0000001110100000,
    64'h0000201111100000,
    64'h0000101211170200,
    64'h0000171221110100,
    64'h0000711211111110,
    64'h0020011111211110,
    64'h0010111211220011,
    64'h0011102211220001,
    64'h0011102201000000,
    64'h0001000000000000,
    64'h0001000000000000,
    // code x02
    64'h0000000000000000,
    64'h0001000000000000,
    64'h0001100000000000,
    64'h0000110000000000,
    64'h0000111102000000,
    64'h0000111117102000,
    64'h0000011111110200,
    64'h0002712211111110,
    64'h0000112111111111,
    64'h0000011111220001,
    64'h0000011111120000,
    64'h0020111211100000,
    64'h0002110220100000,
    64'h0000110000000000,
    64'h0000110000000000,
    64'h0000010000000000,
    // code x03
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0010000000000000,
    64'h0001000020020000,
    64'h0000110001002000,
    64'h0000111007100100,
    64'h0000011111111110,
    64'h0000001221111111,
    64'h0002001211112000,
    64'h0000171111122000,
    64'h0000011111100000,
    64'h0002001112010000,
    64'h0000201122001000,
    64'h0000011100000000,
    64'h0000001100000000,
    64'h0000000100000000,
    // code x04
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000020000,
    64'h0110000200002000,
    64'h0011110710011110,
    64'h0001111111111111,
    64'h0000111221110000,
    64'h0000111211122000,
    64'h0000011111112000,
    64'h0000271111110000,
    64'h0000011112111000,
    64'h0000001112200000,
    64'h0000020110000000,
    64'h0000002110000000,
    64'h0000000110000000,
    64'h0000000011000000,
    // code x05
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000211100,
    64'h0000000000001111,
    64'h0000002117011100,
    64'h0001100071110000,
    64'h1111111111112200,
    64'h0001111222122200,
    64'h0000011121111000,
    64'h0000001111111100,
    64'h0000211111222000,
    64'h0000000711122000,
    64'h0000000001100000,
    64'h0000000211100000,
    64'h0000000001110000,
    64'h0000000000011000,
    // code x06
    64'h0000000022111111,
    64'h0000000000001110,
    64'h0000000000011100,
    64'h0000022117111000,
    64'h0000000071111220,
    64'h0000000111112220,
    64'h0001111112211100,
    64'h1111111122111111,
    64'h0001111112211100,
    64'h0000000111112220,
    64'h0000000071111220,
    64'h0000022117111000,
    64'h0000000000011100,
    64'h0000000000001110,
    64'h0000000022111111,
    64'h0000000000000000,
    // code x07
    64'h0000000200000000,
    64'h0000000200000000,
    64'h0000000200000000,
    64'h0000002220000000,
    64'h0000002220000000,
    64'h0008002220080000,
    64'h0008002220080000,
    64'h0002022222020000,
    64'h8002722822720080,
    64'h8007228882270080,
    64'h2002228282220020,
    64'h2022222222222020,
    64'h2222282228222220,
    64'h2220882228802220,
    64'h2200880208800220,
    64'h2000000200000020,
    // code x08
    64'h0000002000000000,
    64'h0000002000000000,
    64'h0000002000000000,
    64'h0000022200000000,
    64'h0000022200800000,
    64'h0000002220200000,
    64'h0000802222200000,
    64'h0000202822270800,
    64'h0000272882220200,
    64'h0000722822222220,
    64'h0080022222822220,
    64'h0020222822880022,
    64'h0022208822880002,
    64'h0022208802000000,
    64'h0002000000000000,
    64'h0002000000000000,
    // code x09
    64'h0000000000000000,
    64'h0002000000000000,
    64'h0002200000000000,
    64'h0000220000000000,
    64'h0000222208000000,
    64'h0000222227208000,
    64'h0000022222220800,
    64'h0008728822222220,
    64'h0000228222222222,
    64'h0000022222880002,
    64'h0000022222280000,
    64'h0080222822200000,
    64'h0008220880200000,
    64'h0000220000000000,
    64'h0000220000000000,
    64'h0000020000000000,
    // code x0A
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0020000000000000,
    64'h0002000080080000,
    64'h0000220002008000,
    64'h0000222007200200,
    64'h0000022222222220,
    64'h0000002882222222,
    64'h0008002822228000,
    64'h0000272222288000,
    64'h0000022222200000,
    64'h0008002228020000,
    64'h0000802288002000,
    64'h0000022200000000,
    64'h0000002200000000,
    64'h0000000200000000,
    // code x0B
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000080000,
    64'h0220000800008000,
    64'h0022220720022220,
    64'h0002222222222222,
    64'h0000222882220000,
    64'h0000222822288000,
    64'h0000022222228000,
    64'h0000872222220000,
    64'h0000022228222000,
    64'h0000002228800000,
    64'h0000080220000000,
    64'h0000008220000000,
    64'h0000000220000000,
    64'h0000000022000000,
    // code x0C
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000822200,
    64'h0000000000002222,
    64'h0000008227022200,
    64'h0002200072220000,
    64'h2222222222228800,
    64'h0002222888288800,
    64'h0000022282222000,
    64'h0000002222222200,
    64'h0000822222888000,
    64'h0000000722288000,
    64'h0000000002200000,
    64'h0000000822200000,
    64'h0000000002220000,
    64'h0000000000022000,
    // code x0D
    64'h0000000088222222,
    64'h0000000000002220,
    64'h0000000000022200,
    64'h0000088227222000,
    64'h0000000072222880,
    64'h0000000222228880,
    64'h0002222228822200,
    64'h2222222288222222,
    64'h0002222228822200,
    64'h0000000222228880,
    64'h0000000072222880,
    64'h0000088227222000,
    64'h0000000000022200,
    64'h0000000000002220,
    64'h0000000088222222,
    64'h0000000000000000,
    // code x0E
    64'h0000000000000000,
    64'h0000000606000000,
    64'h0000663363366000,
    64'h0000063363360000,
    64'h0000006666600000,
    64'h0000664464466000,
    64'h0006664444466600,
    64'h0666664444466666,
    64'h0066604444406660,
    64'h0006600303006600,
    64'h0006600303006600,
    64'h0006660000066600,
    64'h0000660000066000,
    64'h0000066000660000,
    64'h0000006606600000,
    64'h0000000606000000,
    // code x0F
    64'h0000000606000000,
    64'h0000000606000000,
    64'h0000663363366000,
    64'h0000063363360000,
    64'h0000006666600000,
    64'h0000064464460000,
    64'h0006664444466600,
    64'h0666664444466666,
    64'h0066664444466660,
    64'h0063660303066360,
    64'h0663600303006366,
    64'h0636600000006636,
    64'h0633600000006336,
    64'h0633600000006336,
    64'h0666600000006666,
    64'h0066000000000660,
    // code x10
    64'h0000000000000000,
    64'h0000000600600000,
    64'h0000066336000000,
    64'h0066336330000000,
    64'h0006636666660000,
    64'h0000064644666060,
    64'h0006644444666600,
    64'h0006644444406600,
    64'h0066664444006600,
    64'h0666604303006600,
    64'h0066600303066600,
    64'h0006600000006600,
    64'h0006666000066000,
    64'h0000066600060000,
    64'h0000006660600000,
    64'h0000000060000000,
    // code x11
    64'h0000000000000000,
    64'h0000600600000000,
    64'h0006633600000000,
    64'h0003636006660000,
    64'h0663664466660000,
    64'h0006644446666000,
    64'h0000444446666600,
    64'h0006644430066360,
    64'h0066643030063360,
    64'h0666660000006660,
    64'h0006360000006660,
    64'h0006360000000000,
    64'h0006336000000000,
    64'h0006666000000000,
    64'h0000666000000000,
    64'h0000060000000000,
    // code x12
    64'h0000000000000000,
    64'h0000000600000000,
    64'h0000000600000000,
    64'h0000633006606600,
    64'h0006033666666000,
    64'h0003366446666000,
    64'h0003366444066600,
    64'h0660644444406660,
    64'h0000644444306660,
    64'h0006664440300660,
    64'h0006660433000660,
    64'h0000666000000600,
    64'h0006666660000600,
    64'h0006006666666000,
    64'h0000000666600000,
    64'h0000000000000000,
    // code x13
    64'h0000000000000000,
    64'h0000600006000000,
    64'h0000600066000000,
    64'h0063360666666600,
    64'h0666664666333660,
    64'h0033644446663666,
    64'h0036444430006660,
    64'h0660444400000000,
    64'h0000644330000000,
    64'h0006666000000000,
    64'h0006666000000000,
    64'h0006666660000000,
    64'h0000066636600000,
    64'h0000006336600000,
    64'h0000000666600000,
    64'h0000000000000000,
    // code x14
    64'h0000000000000000,
    64'h0000000006000000,
    64'h0006000066600000,
    64'h0006606666666000,
    64'h0003606666666000,
    64'h0063364460006600,
    64'h0066644444006660,
    64'h0633664443300660,
    64'h0033644440000066,
    64'h0060644443300000,
    64'h0600666400000060,
    64'h0000666000606600,
    64'h0000066666666000,
    64'h0000006666660000,
    64'h0000060000000000,
    64'h0000000000000000,
    // code x15
    64'h0000000000000000,
    64'h0000000600666660,
    64'h0000000666633366,
    64'h0000006663363366,
    64'h0060006666666660,
    64'h0066066666000000,
    64'h0033644440000000,
    64'h6633644443300000,
    64'h0066664440000000,
    64'h6633644443300000,
    64'h0033644440000000,
    64'h0066066666000000,
    64'h0060006666666660,
    64'h0000006663363366,
    64'h0000000666633366,
    64'h0000000600666660,
    // code x16
    64'h0000000000000000,
    64'h0000000707000000,
    64'h000077bb7bb77000,
    64'h000007bb7bb70000,
    64'h0000007777700000,
    64'h000077aa7aa77000,
    64'h000777aaaaa77700,
    64'h077777aaaaa77777,
    64'h007770aaaaa07770,
    64'h0007700b0b007700,
    64'h0007700b0b007700,
    64'h0007770000077700,
    64'h0000770000077000,
    64'h0000077000770000,
    64'h0000007707700000,
    64'h0000000707000000,
    // code x17
    64'h0000000707000000,
    64'h0000000707000000,
    64'h000077bb7bb77000,
    64'h000007bb7bb70000,
    64'h0000007777700000,
    64'h000007aa7aa70000,
    64'h000777aaaaa77700,
    64'h077777aaaaa77777,
    64'h007777aaaaa77770,
    64'h007b770b0b077b70,
    64'h077b700b0b007b77,
    64'h07b77000000077b7,
    64'h07bb700000007bb7,
    64'h07bb700000007bb7,
    64'h0777700000007777,
    64'h0077000000000770,
    // code x18
    64'h0000000000000000,
    64'h0000000700700000,
    64'h0000077bb7000000,
    64'h0077bb7bb0000000,
    64'h00077b7777770000,
    64'h000007a7aa777070,
    64'h00077aaaaa777700,
    64'h00077aaaaaa07700,
    64'h007777aaaa007700,
    64'h077770ab0b007700,
    64'h0077700b0b077700,
    64'h0007700000007700,
    64'h0007777000077000,
    64'h0000077700070000,
    64'h0000007770700000,
    64'h0000000070000000,
    // code x19
    64'h0000000000000000,
    64'h0000700700000000,
    64'h00077bb700000000,
    64'h000b7b7007770000,
    64'h077b77aa77770000,
    64'h00077aaaa7777000,
    64'h0000aaaaa7777700,
    64'h00077aaab0077b70,
    64'h00777ab0b007bb70,
    64'h0777770000007770,
    64'h0007b70000007770,
    64'h0007b70000000000,
    64'h0007bb7000000000,
    64'h0007777000000000,
    64'h0000777000000000,
    64'h0000070000000000,
    // code x1A
    64'h0000000000000000,
    64'h0000000700000000,
    64'h0000000700000000,
    64'h00007bb007707700,
    64'h00070bb777777000,
    64'h000bb77aa7777000,
    64'h000bb77aaa077700,
    64'h07707aaaaaa07770,
    64'h00007aaaaab07770,
    64'h000777aaa0b00770,
    64'h0007770abb000770,
    64'h0000777000000700,
    64'h0007777770000700,
    64'h0007007777777000,
    64'h0000000777700000,
    64'h0000000000000000,
    // code x1B
    64'h0000000000000000,
    64'h0000700007000000,
    64'h0000700077000000,
    64'h007bb70777777700,
    64'h077777a777bbb770,
    64'h00bb7aaaa777b777,
    64'h00b7aaaab0007770,
    64'h0770aaaa00000000,
    64'h00007aabb0000000,
    64'h0007777000000000,
    64'h0007777000000000,
    64'h0007777770000000,
    64'h00000777b7700000,
    64'h0000007bb7700000,
    64'h0000000777700000,
    64'h0000000000000000,
    // code x1C
    64'h0000000000000000,
    64'h0000000007000000,
    64'h0007000077700000,
    64'h0007707777777000,
    64'h000b707777777000,
    64'h007bb7aa70007700,
    64'h00777aaaaa007770,
    64'h07bb77aaabb00770,
    64'h00bb7aaaa0000077,
    64'h00707aaaabb00000,
    64'h0700777a00000070,
    64'h0000777000707700,
    64'h0000077777777000,
    64'h0000007777770000,
    64'h0000070000000000,
    64'h0000000000000000,
    // code x1D
    64'h0000000000000000,
    64'h0000000700777770,
    64'h00000007777bbb77,
    64'h000000777bb7bb77,
    64'h0070007777777770,
    64'h0077077777000000,
    64'h00bb7aaaa0000000,
    64'h77bb7aaaabb00000,
    64'h007777aaa0000000,
    64'h77bb7aaaabb00000,
    64'h00bb7aaaa0000000,
    64'h0077077777000000,
    64'h0070007777777770,
    64'h000000777bb7bb77,
    64'h00000007777bbb77,
    64'h0000000700777770,
    // code x1E
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000200000002000,
    64'h0000200707002000,
    64'h0000201212102000,
    64'h0000201111102000,
    64'h0000222111222000,
    64'h0000002777200000,
    64'h0000222777222000,
    64'h0000222111222000,
    64'h0000220777022000,
    64'h0000220070022000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    // code x1F
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000200707002000,
    64'h0022200707002220,
    64'h0022201212102220,
    64'h0022201111102220,
    64'h0002222111222200,
    64'h0000222777222000,
    64'h0002222777222200,
    64'h0022222111222220,
    64'h0002220777022200,
    64'h0000020000020000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    // code x20
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000200000,
    64'h0000000000200000,
    64'h0020000700200000,
    64'h0020071210020000,
    64'h0020127777220000,
    64'h0002077772000000,
    64'h0002221112220000,
    64'h0000021111220000,
    64'h0000222777222000,
    64'h0000222777022000,
    64'h0000220070000000,
    64'h0000220000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    // code x21
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000002020000,
    64'h0000007002222000,
    64'h0000700700222000,
    64'h0000070210022000,
    64'h0020021112222000,
    64'h0222011112222220,
    64'h0222022177222200,
    64'h0222222771122220,
    64'h0002222211702000,
    64'h0000222217700000,
    64'h0000222200700000,
    64'h0000000200000000,
    64'h0000000000000000,
    64'h0000000000000000,
    // code x22
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000220000000,
    64'h0000000022000000,
    64'h0000070102200000,
    64'h0000702102000000,
    64'h0000021112022000,
    64'h0020111177222200,
    64'h0022001777102200,
    64'h0002222771170000,
    64'h0000200211770000,
    64'h0000002207770000,
    64'h0000002220000000,
    64'h0000000220000000,
    64'h0000000000000000,
    64'h0000000000000000,
    // code x23
    64'h0000000000000000,
    64'h0000000222000000,
    64'h0000002222000000,
    64'h0000000222200000,
    64'h0000700002222000,
    64'h0000072122222000,
    64'h0007001122222000,
    64'h0000721117222200,
    64'h0000011177110000,
    64'h0022002271170000,
    64'h0002202221777000,
    64'h0022222222000000,
    64'h0002222222200000,
    64'h0000000222000000,
    64'h0000000202000000,
    64'h0000000000000000,
    // code x24
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000222000000000,
    64'h0000000220000000,
    64'h0000001020222200,
    64'h0000072722222200,
    64'h0000017711220000,
    64'h0000727711770000,
    64'h0000017711777000,
    64'h0000007221770000,
    64'h0022202022200000,
    64'h0000022022220000,
    64'h0000000000220000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    // code x25
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000222000200000,
    64'h0000222202220000,
    64'h0002222222220000,
    64'h0000000222222000,
    64'h0000011222200000,
    64'h0007721177170000,
    64'h0000011177170000,
    64'h0007721177170000,
    64'h0000011222200000,
    64'h0000000222222000,
    64'h0002222222220000,
    64'h0000222202220000,
    64'h0000222000200000,
    64'h0000000000000000,
    // code x26
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000700040007000,
    64'h0000704242407000,
    64'h0000072242270000,
    64'h0000004444400000,
    64'h0000077444770000,
    64'h0000077222770000,
    64'h0000770222077000,
    64'h0000770444077000,
    64'h0000770222077000,
    64'h0000770020077000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    // code x27
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0007000040000700,
    64'h0000704242407000,
    64'h0000072242270000,
    64'h0000004444400000,
    64'h0000077444770000,
    64'h0000777222777000,
    64'h0007770222077700,
    64'h0077770444077770,
    64'h0077700222007770,
    64'h0077700020007770,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    // code x28
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000070000,
    64'h0000000400070000,
    64'h0000002424700000,
    64'h0007042422000000,
    64'h0000774444770000,
    64'h0000004444770000,
    64'h0000077222077000,
    64'h0000077222207700,
    64'h0000077044407700,
    64'h0000077022207700,
    64'h0000077002000000,
    64'h0000077000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    // code x29
    64'h0000000000000000,
    64'h0000000007000000,
    64'h0000040407000000,
    64'h0000042270000000,
    64'h0000424447000000,
    64'h0770224447777700,
    64'h0007044427777770,
    64'h0000772222077770,
    64'h0000777244000770,
    64'h0000770442200000,
    64'h0000777022000000,
    64'h0007770000000000,
    64'h0007777000000000,
    64'h0000770000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    // code x2A
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000700000000,
    64'h0000000070000000,
    64'h0000402470000000,
    64'h0000042247000000,
    64'h0000224447777000,
    64'h0070424442477700,
    64'h0007744422477770,
    64'h0000077224420700,
    64'h0000007444200000,
    64'h0000007772020000,
    64'h0000007770000000,
    64'h0000000777000000,
    64'h0000000070000000,
    64'h0000000000000000,
    // code x2B
    64'h0000000000000000,
    64'h0000070000000000,
    64'h0000070000000000,
    64'h0000007000077000,
    64'h0000420777777700,
    64'h0044224777777700,
    64'h0002444270707000,
    64'h0042444224000000,
    64'h0007442244200000,
    64'h0770777242200000,
    64'h0000077002000000,
    64'h0000077700000000,
    64'h0000077700000000,
    64'h0000077770000000,
    64'h0000007770000000,
    64'h0000000000000000,
    // code x2C
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000070000000000,
    64'h0000007000000000,
    64'h0000047077777700,
    64'h0000224477777700,
    64'h0004444422000000,
    64'h0000224422420000,
    64'h0000424422422000,
    64'h0000707702420000,
    64'h0077007770000000,
    64'h0000000077770000,
    64'h0000000007770000,
    64'h0000000000000000,
    64'h0000000000000000,
    // code x2D
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000777000,
    64'h0007000007777000,
    64'h0000700077777000,
    64'h0000070777700000,
    64'h0000424770000000,
    64'h0000224422420000,
    64'h0004444422422000,
    64'h0000224422420000,
    64'h0000424770000000,
    64'h0000070777700000,
    64'h0000700077777000,
    64'h0007000007777000,
    64'h0000000000777000,
    64'h0000000000000000,
    // code x2E
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000700000000,
    64'h0000000700000000,
    64'h0000007770000000,
    64'h0000007170000000,
    64'h0000000200000000,
    64'h0000000200000000,
    64'h0000000200000000,
    64'h0000000200000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    // code x2F
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000100000000,
    64'h0000000100000000,
    64'h0000000100000000,
    64'h0000000100000000,
    64'h0000002520000000,
    64'h0000002220000000,
    64'h0000000200000000,
    64'h0000000200000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    // code x30
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000200000000,
    64'h0000000200000000,
    64'h0000000200000000,
    64'h0000000200000000,
    64'h0000007170000000,
    64'h0000007770000000,
    64'h0000000700000000,
    64'h0000000700000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    // code x31
    64'h0000000000000000,
    64'h0000000100000000,
    64'h0000000100000000,
    64'h0000001110000000,
    64'h0000001110000000,
    64'h0002001110020000,
    64'h0002001110020000,
    64'h0201011211010200,
    64'h0201712221710200,
    64'h0107112121170100,
    64'h0101111111110100,
    64'h0111121112111100,
    64'h0111221112211100,
    64'h0110220102201100,
    64'h0100000100000100,
    64'h0000000000000000,
    // code x32
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h1111111000000000,
    64'h2222222000000000,
    64'h2222222000000000,
    64'h1111111000000000,
    64'h2222222000000000,
    64'h2222222000000000,
    64'h1111111000000000,
    64'h1911191000000000,
    64'h1191911000000000,
    64'h0119110000000000,
    64'h0011100000000000,
    64'h0001000000000000
  };

  assign data_o = ROM[addr_i];

endmodule
