module font_rom (
  input [7:0] addr_i,
  output [7:0] data_o
);

localparam int AddrWidth = 8;
localparam int DataWidth = 8;

localparam logic [0:2**AddrWidth-1][DataWidth-1:0] ROM = {
  // code x00
  8'b00000000, // 0
  8'b00000000, // 1
  8'b01111100, // 2  *****
  8'b11000110, // 3 **   **
  8'b11000110, // 4 **   **
  8'b01100000, // 5  **
  8'b00111000, // 6   ***
  8'b00001100, // 7     **
  8'b00000110, // 8      **
  8'b11000110, // 9 **   **
  8'b11000110, // a **   **
  8'b01111100, // b  *****
  8'b00000000, // c
  8'b00000000, // d
  8'b00000000, // e
  8'b00000000, // f
  // code x01
  8'b00000000, // 0
  8'b00000000, // 1
  8'b00111100, // 2   ****
  8'b01100110, // 3  **  **
  8'b11000010, // 4 **    *
  8'b11000000, // 5 **
  8'b11000000, // 6 **
  8'b11000000, // 7 **
  8'b11000000, // 8 **
  8'b11000010, // 9 **    *
  8'b01100110, // a  **  **
  8'b00111100, // b   ****
  8'b00000000, // c
  8'b00000000, // d
  8'b00000000, // e
  8'b00000000, // f
  // code x02
  8'b00000000, // 0
  8'b00000000, // 1
  8'b01111100, // 2  *****
  8'b11000110, // 3 **   **
  8'b11000110, // 4 **   **
  8'b11000110, // 5 **   **
  8'b11000110, // 6 **   **
  8'b11000110, // 7 **   **
  8'b11000110, // 8 **   **
  8'b11000110, // 9 **   **
  8'b11000110, // a **   **
  8'b01111100, // b  *****
  8'b00000000, // c
  8'b00000000, // d
  8'b00000000, // e
  8'b00000000, // f
  // code x03
  8'b00000000, // 0
  8'b00000000, // 1
  8'b11111100, // 2 ******
  8'b01100110, // 3  **  **
  8'b01100110, // 4  **  **
  8'b01100110, // 5  **  **
  8'b01111100, // 6  *****
  8'b01101100, // 7  ** **
  8'b01100110, // 8  **  **
  8'b01100110, // 9  **  **
  8'b01100110, // a  **  **
  8'b11100110, // b ***  **
  8'b00000000, // c
  8'b00000000, // d
  8'b00000000, // e
  8'b00000000, // f
  // code x04
  8'b00000000, // 0
  8'b00000000, // 1
  8'b11111110, // 2 *******
  8'b01100110, // 3  **  **
  8'b01100010, // 4  **   *
  8'b01101000, // 5  ** *
  8'b01111000, // 6  ****
  8'b01101000, // 7  ** *
  8'b01100000, // 8  **
  8'b01100010, // 9  **   *
  8'b01100110, // a  **  **
  8'b11111110, // b *******
  8'b00000000, // c
  8'b00000000, // d
  8'b00000000, // e
  8'b00000000, // f
  // code x05
  8'b00000000, // 0
  8'b00000000, // 1
  8'b00000000, // 2
  8'b00000000, // 3
  8'b00011000, // 4    **
  8'b00011000, // 5    **
  8'b00000000, // 6
  8'b00000000, // 7
  8'b00000000, // 8
  8'b00011000, // 9    **
  8'b00011000, // a    **
  8'b00000000, // b
  8'b00000000, // c
  8'b00000000, // d
  8'b00000000, // e
  8'b00000000, // f
  // code x06
  8'b00000000, // 0
  8'b00000000, // 1
  8'b01111100, // 2  *****
  8'b11000110, // 3 **   **
  8'b11000110, // 4 **   **
  8'b11001110, // 5 **  ***
  8'b11011110, // 6 ** ****
  8'b11110110, // 7 **** **
  8'b11100110, // 8 ***  **
  8'b11000110, // 9 **   **
  8'b11000110, // a **   **
  8'b01111100, // b  *****
  8'b00000000, // c
  8'b00000000, // d
  8'b00000000, // e
  8'b00000000, // f
  // code x07
  8'b00000000, // 0
  8'b00000000, // 1
  8'b00011000, // 2
  8'b00111000, // 3
  8'b01111000, // 4    **
  8'b00011000, // 5   ***
  8'b00011000, // 6  ****
  8'b00011000, // 7    **
  8'b00011000, // 8    **
  8'b00011000, // 9    **
  8'b00011000, // a    **
  8'b01111110, // b    **
  8'b00000000, // c    **
  8'b00000000, // d  ******
  8'b00000000, // e
  8'b00000000, // f
  // code x08
  8'b00000000, // 0
  8'b00000000, // 1
  8'b01111100, // 2  *****
  8'b11000110, // 3 **   **
  8'b00000110, // 4      **
  8'b00001100, // 5     **
  8'b00011000, // 6    **
  8'b00110000, // 7   **
  8'b01100000, // 8  **
  8'b11000000, // 9 **
  8'b11000110, // a **   **
  8'b11111110, // b *******
  8'b00000000, // c
  8'b00000000, // d
  8'b00000000, // e
  8'b00000000, // f
  // code x09
  8'b00000000, // 0
  8'b00000000, // 1
  8'b01111100, // 2  *****
  8'b11000110, // 3 **   **
  8'b00000110, // 4      **
  8'b00000110, // 5      **
  8'b00111100, // 6   ****
  8'b00000110, // 7      **
  8'b00000110, // 8      **
  8'b00000110, // 9      **
  8'b11000110, // a **   **
  8'b01111100, // b  *****
  8'b00000000, // c
  8'b00000000, // d
  8'b00000000, // e
  8'b00000000, // f
  // code x0A
  8'b00000000, // 0
  8'b00000000, // 1
  8'b00001100, // 2     **
  8'b00011100, // 3    ***
  8'b00111100, // 4   ****
  8'b01101100, // 5  ** **
  8'b11001100, // 6 **  **
  8'b11111110, // 7 *******
  8'b00001100, // 8     **
  8'b00001100, // 9     **
  8'b00001100, // a     **
  8'b00011110, // b    ****
  8'b00000000, // c
  8'b00000000, // d
  8'b00000000, // e
  8'b00000000, // f
  // code x0B
  8'b00000000, // 0
  8'b00000000, // 1
  8'b11111110, // 2 *******
  8'b11000000, // 3 **
  8'b11000000, // 4 **
  8'b11000000, // 5 **
  8'b11111100, // 6 ******
  8'b00000110, // 7      **
  8'b00000110, // 8      **
  8'b00000110, // 9      **
  8'b11000110, // a **   **
  8'b01111100, // b  *****
  8'b00000000, // c
  8'b00000000, // d
  8'b00000000, // e
  8'b00000000, // f
  // code x0C
  8'b00000000, // 0
  8'b00000000, // 1
  8'b00111000, // 2   ***
  8'b01100000, // 3  **
  8'b11000000, // 4 **
  8'b11000000, // 5 **
  8'b11111100, // 6 ******
  8'b11000110, // 7 **   **
  8'b11000110, // 8 **   **
  8'b11000110, // 9 **   **
  8'b11000110, // a **   **
  8'b01111100, // b  *****
  8'b00000000, // c
  8'b00000000, // d
  8'b00000000, // e
  8'b00000000, // f
  // code x0D
  8'b00000000, // 0
  8'b00000000, // 1
  8'b11111110, // 2 *******
  8'b11000110, // 3 **   **
  8'b00000110, // 4      **
  8'b00000110, // 5      **
  8'b00001100, // 6     **
  8'b00011000, // 7    **
  8'b00110000, // 8   **
  8'b00110000, // 9   **
  8'b00110000, // a   **
  8'b00110000, // b   **
  8'b00000000, // c
  8'b00000000, // d
  8'b00000000, // e
  8'b00000000, // f
  // code x0E
  8'b00000000, // 0
  8'b00000000, // 1
  8'b01111100, // 2  *****
  8'b11000110, // 3 **   **
  8'b11000110, // 4 **   **
  8'b11000110, // 5 **   **
  8'b01111100, // 6  *****
  8'b11000110, // 7 **   **
  8'b11000110, // 8 **   **
  8'b11000110, // 9 **   **
  8'b11000110, // a **   **
  8'b01111100, // b  *****
  8'b00000000, // c
  8'b00000000, // d
  8'b00000000, // e
  8'b00000000, // f
  // code x0F
  8'b00000000, // 0
  8'b00000000, // 1
  8'b01111100, // 2  *****
  8'b11000110, // 3 **   **
  8'b11000110, // 4 **   **
  8'b11000110, // 5 **   **
  8'b01111110, // 6  ******
  8'b00000110, // 7      **
  8'b00000110, // 8      **
  8'b00000110, // 9      **
  8'b00001100, // a     **
  8'b01111000, // b  ****
  8'b00000000, // c
  8'b00000000, // d
  8'b00000000, // e
  8'b00000000  // f
};

assign data_o = ROM[addr_i];

endmodule
